`timescale 1ns / 1ps

module fpga_ip_example_tb();
endmodule
