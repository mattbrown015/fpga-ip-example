`timescale 1ns / 1ps

module fpga_ip_example(
    input clk_in1_p,
    input clk_in1_n
    );
endmodule
